-- Copyright (C) 2017  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Intel and sold by Intel or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- Generated by Quartus Prime Version 17.0.0 Build 595 04/25/2017 SJ Lite Edition
-- Created on Mon Oct  9 17:52:23 2017

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY CronoSM IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        ent : IN STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
        buttons : IN STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
        mux : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
        enable : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
        rst : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
    );
END CronoSM;

ARCHITECTURE BEHAVIOR OF CronoSM IS
    TYPE type_fstate IS (state1,state2,state3,state4,state5,state6,state7,state0,stateZerar);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,ent,buttons)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state0;
            mux <= "000";
            enable <= "000000";
            rst <= "000000";
        ELSE
            mux <= "000";
            enable <= "000000";
            rst <= "000000";
            CASE fstate IS
                WHEN state1 =>
                    IF (((ent(3 DOWNTO 0) = "1001") AND (buttons(1 DOWNTO 0) /= "01"))) THEN
                        reg_fstate <= state2;
                    ELSIF ((buttons(1 DOWNTO 0) = "01")) THEN
                        reg_fstate <= state0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    mux <= "000";

                    enable <= "000001";

                    rst <= "000000";
                WHEN state2 =>
                    IF ((ent(3 DOWNTO 0) = "0110")) THEN
                        reg_fstate <= state3;
                    ELSIF ((ent(3 DOWNTO 0) < "0110")) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    mux <= "001";

                    enable <= "000010";

                    rst <= "000001";
                WHEN state3 =>
                    IF ((ent(3 DOWNTO 0) = "1010")) THEN
                        reg_fstate <= state4;
                    ELSIF ((ent(3 DOWNTO 0) < "1010")) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    mux <= "010";

                    enable <= "000100";

                    rst <= "000010";
                WHEN state4 =>
                    IF ((ent(3 DOWNTO 0) = "0110")) THEN
                        reg_fstate <= state5;
                    ELSIF ((ent(3 DOWNTO 0) < "0110")) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state4;
                    END IF;

                    mux <= "011";

                    enable <= "001000";

                    rst <= "000100";
                WHEN state5 =>
                    IF ((ent(3 DOWNTO 0) = "1010")) THEN
                        reg_fstate <= state6;
                    ELSIF ((ent(3 DOWNTO 0) < "1010")) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state5;
                    END IF;

                    mux <= "100";

                    enable <= "010000";

                    rst <= "001000";
                WHEN state6 =>
                    IF ((ent(3 DOWNTO 0) < "0010")) THEN
                        reg_fstate <= state1;
                    ELSIF ((ent(3 DOWNTO 0) = "0010")) THEN
                        reg_fstate <= state7;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state6;
                    END IF;

                    mux <= "101";

                    enable <= "100000";

                    rst <= "010000";
                WHEN state7 =>
                    reg_fstate <= state1;

                    mux <= "000";

                    enable <= "000000";

                    rst <= "100000";
                WHEN state0 =>
                    IF ((buttons(1 DOWNTO 0) = "10")) THEN
                        reg_fstate <= stateZerar;
                    ELSIF ((buttons(1 DOWNTO 0) = "01")) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state0;
                    END IF;
                WHEN stateZerar =>
                    reg_fstate <= state0;

                    rst <= "111111";
                WHEN OTHERS => 
                    mux <= "XXX";
                    enable <= "XXXXXX";
                    rst <= "XXXXXX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
