-- Copyright (C) 2017  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Intel and sold by Intel or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- Generated by Quartus Prime Version 17.0.0 Build 595 04/25/2017 SJ Lite Edition
-- Created on Sun Oct  8 19:40:05 2017

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ModoSM IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        ajusteMux : IN STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
        ajusteEnable : IN STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
        ajusteRst : IN STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
        ajuste : IN STD_LOGIC := '0';
        relEnable : IN STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
        relMux : IN STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
        relRst : IN STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
        ajusteClock : IN STD_LOGIC := '0';
        relClock : IN STD_LOGIC := '0';
        muxout : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
        enableout : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
        rstout : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
        clockOut : OUT STD_LOGIC
    );
END ModoSM;

ARCHITECTURE BEHAVIOR OF ModoSM IS
    TYPE type_fstate IS (state1,state2);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,ajusteMux,ajusteEnable,ajusteRst,ajuste,relEnable,relMux,relRst,ajusteClock,relClock)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            muxout <= "000";
            enableout <= "000000";
            rstout <= "000000";
            clockOut <= '0';
        ELSE
            muxout <= "000";
            enableout <= "000000";
            rstout <= "000000";
            clockOut <= '0';
            CASE fstate IS
                WHEN state1 =>
                    IF ((ajuste = '1')) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    enableout <= relEnable(5 DOWNTO 0);

                    muxout <= relMux(2 DOWNTO 0);

                    rstout <= relRst(5 DOWNTO 0);

                    clockOut <= relClock;
                WHEN state2 =>
                    IF (NOT((ajuste = '1'))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    enableout <= ajusteEnable(5 DOWNTO 0);

                    muxout <= ajusteMux(2 DOWNTO 0);

                    rstout <= ajusteRst(5 DOWNTO 0);

                    clockOut <= ajusteClock;
                WHEN OTHERS => 
                    muxout <= "XXX";
                    enableout <= "XXXXXX";
                    rstout <= "XXXXXX";
                    clockOut <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
