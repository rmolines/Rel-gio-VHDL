-- Copyright (C) 2017  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Intel and sold by Intel or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- Generated by Quartus Prime Version 17.0.0 Build 595 04/25/2017 SJ Lite Edition
-- Created on Mon Oct  9 18:01:47 2017

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY AlarmeSM IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        a : IN STD_LOGIC_VECTOR(23 DOWNTO 0) := "000000000000000000000000";
        b : IN STD_LOGIC_VECTOR(23 DOWNTO 0) := "000000000000000000000000";
        estado : IN STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
        c : IN STD_LOGIC_VECTOR(23 DOWNTO 0) := "000000000000000000000000";
        d : OUT STD_LOGIC_VECTOR(23 DOWNTO 0)
    );
END AlarmeSM;

ARCHITECTURE BEHAVIOR OF AlarmeSM IS
    TYPE type_fstate IS (state1,state2,state3);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,a,b,estado,c)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            d <= "000000000000000000000000";
        ELSE
            d <= "000000000000000000000000";
            CASE fstate IS
                WHEN state1 =>
                    IF ((estado(1 DOWNTO 0) = "01")) THEN
                        reg_fstate <= state2;
                    ELSIF ((estado(1 DOWNTO 0) = "10")) THEN
                        reg_fstate <= state3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    d <= a(23 DOWNTO 0);
                WHEN state2 =>
                    IF ((estado(1 DOWNTO 0) = "00")) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    d <= b(23 DOWNTO 0);
                WHEN state3 =>
                    IF ((estado(1 DOWNTO 0) = "00")) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    d <= c(23 DOWNTO 0);
                WHEN OTHERS => 
                    d <= "XXXXXXXXXXXXXXXXXXXXXXXX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
